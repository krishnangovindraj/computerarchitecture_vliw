module pipleline_IF_ID( input clk, input reset, input regWrite, input [31:0] instr2Word, output [15:0] p1_aluInstr, output [15:0] p1_memInstr );
	register16bit reg_aluInstr(clk, reset, regWrite, instr2Word[15:0], p1_aluInstr);
	register16bit reg_memInstr(clk, reset, regWrite, instr2Word[31:16], p1_memInstr);
endmodule

module pipeline_ID_EX( 
		input clk, input reset, input regWrite, 
		input [2:0] alu_rn, alu_rm, alu_rd, mem_rn, mem_rd,
		output [2:0] p2_alu_rn, p2_alu_rm, p2_alu_rd, p2_mem_rn, p2_mem_rd,
		
		input [31:0] alu_reg_rm, alu_reg_rn, mem_reg_rn, mem_reg_rd, 
		output [31:0] p2_alu_reg_rm, p2_alu_reg_rns, p2_mem_reg_rn, p2_mem_reg_rd, 
		
		input [31:0] alu_sextImm3, mem_sextImm5, mem_sextImm8,
		output [31:0] p2_alu_sextImm3, p2_mem_sextImm5, p2_mem_sextImm8
	);
	
	register3bit reg_alu_rn( clk, reset, regWrite, 1'b1, alu_rn, p2_alu_rn );
	register3bit reg_alu_rm( clk, reset, regWrite, 1'b1, alu_rm, p2_alu_rm );
	register3bit reg_alu_rd( clk, reset, regWrite, 1'b1, alu_rd, p2_alu_rd );
	
	register3bit reg_mem_rn( clk, reset, regWrite, 1'b1, mem_rn, p2_mem_rn );
	register3bit reg_mem_rd( clk, reset, regWrite, 1'b1, mem_rd, p2_mem_rd );
	
	
	register32bit reg_alu_reg_rn( clk, reset, regWrite, 1'b1, alu_reg_rn, p2_alu_reg_rn );
	register32bit reg_alu_reg_rm( clk, reset, regWrite, 1'b1, alu_reg_rm, p2_alu_reg_rm );
	
	register32bit reg_mem_reg_rn( clk, reset, regWrite, 1'b1, mem_reg_rn, p2_mem_reg_rn );
	register32bit reg_mem_reg_rn( clk, reset, regWrite, 1'b1, mem_reg_rd, p2_mem_reg_rd );
	
	
	register32bit reg_alu_sextImm3( clk, reset, regWrite, 1'b1, alu_sextImm3, p2_alu_sextImm3 );
	register32bit reg_mem_sextImm5( clk, reset, regWrite, 1'b1, mem_sextImm5, p2_mem_sextImm5 );
	register32bit reg_mem_sextImm8( clk, reset, regWrite, 1'b1, mem_sextImm8, p2_mem_sextImm8 );
	
endmodule



